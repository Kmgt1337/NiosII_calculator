library ieee;
use ieee.std_logic_1164.all;

entity seven_segments_contrl_tb is
end entity;

architecture simulation of seven_segments_contrl_tb is

component seven_segments_contrl is
	port
	(
		clk 			: in std_logic;
		neg_in_ena 		: in std_logic;
		neg_ena			: in std_logic;
		number			: in std_logic_vector(10 downto 0);
		
		hex0			: out std_logic_vector(7 downto 0);
		hex1			: out std_logic_vector(7 downto 0);
		hex2			: out std_logic_vector(7 downto 0);
		hex3			: out std_logic_vector(7 downto 0);
		hex4			: out std_logic_vector(7 downto 0);
		hex5			: out std_logic_vector(7 downto 0)
	);
end component;

signal clk : std_logic := '0';
signal neg_in_ena, neg_ena : std_logic;
signal number : std_logic_vector(10 downto 0);
signal hex0, hex1, hex2, hex3, hex4, hex5 : std_logic_vector(7 downto 0);

begin
	uut : seven_segments_contrl 
	port map(clk, neg_in_ena, neg_ena, number, hex0, hex1, hex2, hex3, hex4, hex5);

	clk <= not clk after 1 ns;

	process
	begin
		neg_in_ena <= '0';
		neg_ena <= '0';
		wait for 5 ns;

		number <= "00000000001";
		wait for 5 ns;

		number <= "00000001100";
		wait for 5 ns;

		number <= "00001111011";
		wait for 5 ns;

		number <= "01111111111";
		wait for 5 ns;

		number <= "11111111111";
		neg_ena <= '1';
		wait for 5 ns;

		neg_ena <= '0';
		neg_in_ena <= '1';
		wait for 5 ns;

		neg_ena <= '0';
		neg_in_ena <= '0';
		wait for 200 ns;
	end process;

end architecture;
