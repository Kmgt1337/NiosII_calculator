library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity seven_segments_contrl is
	port
	(
		clk 			: in std_logic;
		neg_in_ena 		: in std_logic;
		neg_ena			: in std_logic;
		number			: in std_logic_vector(10 downto 0);
		
		hex0			: out std_logic_vector(7 downto 0);
		hex1			: out std_logic_vector(7 downto 0);
		hex2			: out std_logic_vector(7 downto 0);
		hex3			: out std_logic_vector(7 downto 0);
		hex4			: out std_logic_vector(7 downto 0);
		hex5			: out std_logic_vector(7 downto 0)
	);
end entity;

architecture behavior of seven_segments_contrl is

component seven_seg is
	port
	(
		neg_ena			: std_logic;
		neg_in_ena		: std_logic;
		inputBCD  		: in std_logic_vector(3 downto 0); -- 4 bits input
		outputHEX 		: out std_logic_vector(7 downto 0) -- 8 bits output
	);
end component;

signal bcd0, bcd1, bcd2, bcd3, bcd4, bcd5 : unsigned(10 downto 0);
signal num_temp : unsigned(10 downto 0);

begin
	process(clk)
	begin
		num_temp <= unsigned(number);
		bcd0 <= num_temp mod 10;
		bcd1 <= (num_temp / 10) mod 10;
		bcd2 <= (num_temp / 100) mod 10;
		bcd3 <= (num_temp / 1000) mod 1000;
	end process;
			
	segment0 : seven_seg 
	port map
	(
		neg_ena => '0',
		neg_in_ena => '0',
		inputBCD => std_logic_vector(bcd0(3 downto 0)),
		outputHEX => hex0
	);

	segment1 : seven_seg 
	port map
	(
		neg_ena => '0',
		neg_in_ena => '0',
		inputBCD => std_logic_vector(bcd1(3 downto 0)),
		outputHEX => hex1
	);

	segment2 : seven_seg 
	port map
	(
		neg_ena => '0',
		neg_in_ena => '0',
		inputBCD => std_logic_vector(bcd2(3 downto 0)),
		outputHEX => hex2
	);

	segment3 : seven_seg 
	port map
	(
		neg_ena => '0',
		neg_in_ena => '0',
		inputBCD => std_logic_vector(bcd3(3 downto 0)),
		outputHEX => hex3
	);

	segment4 : seven_seg 
	port map
	(
		neg_ena => neg_ena,
		neg_in_ena => '0',
		inputBCD => (others => '0'),
		outputHEX => hex4
	);

	segment5 : seven_seg 
	port map
	(
		neg_ena => '0',
		neg_in_ena => neg_in_ena,
		inputBCD => (others => '0'),
		outputHEX => hex5
	);
	
end architecture;