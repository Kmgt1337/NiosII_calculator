
module nios2 (
	clk_clk,
	input_export,
	output_export,
	reset_reset_n);	

	input		clk_clk;
	input	[10:0]	input_export;
	output	[10:0]	output_export;
	input		reset_reset_n;
endmodule
